* NGSPICE file created from ef_smsdac8_ladder.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p35_CN8CXG a_1708_1984# a_712_1984# a_n948_1984#
+ a_n1778_n2416# a_n948_n2416# a_n1446_1984# a_546_1984# a_380_n2416# a_1542_n2416#
+ a_712_n2416# a_n1280_n2416# a_2040_n2416# a_1210_1984# a_n1612_n2416# a_1044_n2416#
+ a_n450_n2416# a_n1944_1984# a_214_n2416# a_n450_1984# a_1044_1984# a_n1778_1984#
+ a_n2110_n2416# a_n284_1984# a_n1114_n2416# a_878_1984# a_1874_n2416# a_2040_1984#
+ a_48_n2416# a_n118_1984# a_1542_1984# a_n1944_n2416# a_1376_n2416# a_n782_n2416#
+ a_n782_1984# a_546_n2416# a_n1280_1984# a_1708_n2416# a_1376_1984# a_380_1984# a_n1446_n2416#
+ a_n2240_n2546# a_n284_n2416# a_n616_1984# a_n616_n2416# a_n1114_1984# a_214_1984#
+ a_1874_1984# a_1210_n2416# a_878_n2416# a_n118_n2416# a_n2110_1984# a_48_1984# a_n1612_1984#
X0 a_n450_1984# a_n450_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X1 a_n1612_1984# a_n1612_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X2 a_n284_1984# a_n284_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X3 a_48_1984# a_48_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X4 a_n948_1984# a_n948_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X5 a_n782_1984# a_n782_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X6 a_1376_1984# a_1376_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X7 a_878_1984# a_878_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X8 a_n1446_1984# a_n1446_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X9 a_n2110_1984# a_n2110_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X10 a_1874_1984# a_1874_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X11 a_n1944_1984# a_n1944_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X12 a_214_1984# a_214_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X13 a_n1280_1984# a_n1280_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X14 a_1210_1984# a_1210_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X15 a_712_1984# a_712_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X16 a_n118_1984# a_n118_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X17 a_n1778_1984# a_n1778_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X18 a_n616_1984# a_n616_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X19 a_1044_1984# a_1044_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X20 a_380_1984# a_380_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X21 a_546_1984# a_546_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X22 a_n1114_1984# a_n1114_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X23 a_1542_1984# a_1542_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X24 a_1708_1984# a_1708_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
X25 a_2040_1984# a_2040_n2416# a_n2240_n2546# sky130_fd_pr__res_high_po_0p35 l=20
.ends

*.subckt ef_smsdac8_ladder
.subckt ef_smsdac8_ladder vdac vdd gnd i_x4[1] i_x1[1] i_x4[0] i_x2[0] i_x2[1] i_x8[0] i_x1[0] i_x8[1]
Xsky130_fd_pr__res_high_po_0p35_CN8CXG_0 vdac m1_2648_n4006# m1_988_610# gnd m1_1652_n4006#
+ m1_988_610# m1_2648_n4006# m1_2648_n4006# i_x1[1] i_x2[0] i_x8[0] gnd m1_2648_n4006#
+ vdd vdac i_x4[1] gnd m1_2648_n4006# m1_1652_n4006# m1_2648_n4006# m1_988_610# gnd
+ m1_1652_n4006# m1_1652_n4006# m1_2648_n4006# gnd gnd m1_2648_n4006# m1_1652_n4006#
+ vdac gnd vdac m1_1652_n4006# m1_988_610# i_x2[1] m1_988_610# i_x1[0] m1_2648_n4006#
+ m1_1652_n4006# i_x8[1] gnd i_x4[0] m1_988_610# m1_1652_n4006# m1_988_610# m1_1652_n4006#
+ gnd vdac vdac m1_2648_n4006# gnd m1_1652_n4006# m1_988_610# sky130_fd_pr__res_high_po_0p35_CN8CXG
.ends

