** sch_path: /home/ejf/Dropbox/Projects/Research_OSIC/TT/tt07-ef-smsdac8-analog/xschem/ef_smsdac8_ladder.sch
.subckt ef_smsdac8_ladder vdac vdd gnd i_x4[1] i_x1[1] i_x4[0] i_x2[0] i_x2[1] i_x8[0] i_x1[0] i_x8[1]
*.PININFO vdd:B vdac:O i_x8[1]:I gnd:B i_x8[0]:I i_x4[1]:I i_x4[0]:I i_x2[1]:I i_x2[0]:I i_x1[1]:I i_x1[0]:I
XR1 i_x8[1] net1 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR6 i_x8[0] net1 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR11 net2 net1 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=4 m=4
XR12 gnd net1 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR16 vdd net1 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR5 i_x4[1] net2 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR22 i_x4[0] net2 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR26 net3 net2 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=4 m=4
XR27 i_x2[1] net3 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR31 i_x2[0] net3 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR35 vdac net3 gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=4 m=4
XR36 i_x1[1] vdac gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR40 i_x1[0] vdac gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR2 gnd gnd gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=2 m=2
XR3 gnd gnd gnd sky130_fd_pr__res_high_po_0p35 L=20 mult=2 m=2
.ends
.end
