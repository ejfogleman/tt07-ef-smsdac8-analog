magic
tech sky130A
magscale 1 2
timestamp 1716599306
<< viali >>
rect 526 668 560 826
rect 4972 668 5006 826
rect 526 -4006 560 -3848
rect 988 -4006 1058 -3574
rect 1154 -4008 1224 -3574
rect 1320 -4006 1390 -3572
rect 1486 -4006 1556 -3572
rect 2316 -4006 2386 -3572
rect 2482 -4006 2552 -3572
rect 3312 -4006 3382 -3572
rect 3478 -4006 3548 -3572
rect 4308 -4006 4378 -3572
rect 4474 -4006 4544 -3572
rect 4972 -4006 5006 -3848
<< metal1 >>
rect 520 826 566 838
rect 4966 826 5012 838
rect 520 668 526 826
rect 560 756 892 826
rect 560 668 566 756
rect 520 656 566 668
rect 988 610 2220 826
rect 2316 610 2398 826
rect 2468 610 3216 826
rect 3312 610 3396 826
rect 3466 610 4212 826
rect 4308 610 4392 826
rect 4462 610 4544 826
rect 4640 756 4972 826
rect 4966 668 4972 756
rect 5006 668 5012 826
rect 4966 656 5012 668
rect 982 -3574 1064 -3562
rect 1148 -3574 1230 -3562
rect 1314 -3572 1396 -3560
rect 1480 -3572 1562 -3560
rect 2310 -3572 2392 -3560
rect 2476 -3572 2558 -3560
rect 3306 -3572 3388 -3560
rect 3472 -3572 3554 -3560
rect 4302 -3572 4384 -3560
rect 4468 -3572 4550 -3560
rect 520 -3848 566 -3836
rect 520 -4006 526 -3848
rect 560 -3936 566 -3848
rect 978 -3936 988 -3574
rect 560 -4006 988 -3936
rect 1058 -4006 1068 -3574
rect 520 -4018 566 -4006
rect 982 -4018 1064 -4006
rect 1144 -4008 1154 -3574
rect 1224 -4008 1234 -3574
rect 1310 -4006 1320 -3572
rect 1390 -4006 1400 -3572
rect 1476 -4006 1486 -3572
rect 1556 -4006 1566 -3572
rect 1652 -4006 1902 -3790
rect 1972 -4006 2220 -3790
rect 2306 -4006 2316 -3572
rect 2386 -4006 2396 -3572
rect 2472 -4006 2482 -3572
rect 2552 -4006 2562 -3572
rect 2648 -4006 2896 -3790
rect 2966 -4006 3216 -3790
rect 3302 -4006 3312 -3572
rect 3382 -4006 3392 -3572
rect 3468 -4006 3478 -3572
rect 3548 -4006 3558 -3572
rect 3644 -4006 3892 -3790
rect 3962 -4006 4212 -3790
rect 4298 -4006 4308 -3572
rect 4378 -4006 4388 -3572
rect 4464 -4006 4474 -3572
rect 4544 -4006 4554 -3572
rect 4966 -3848 5012 -3836
rect 4966 -3936 4972 -3848
rect 4640 -4006 4972 -3936
rect 5006 -4006 5012 -3848
rect 1148 -4020 1230 -4008
rect 1314 -4018 1396 -4006
rect 1480 -4018 1562 -4006
rect 2310 -4018 2392 -4006
rect 2476 -4018 2558 -4006
rect 3306 -4018 3388 -4006
rect 3472 -4018 3554 -4006
rect 4302 -4018 4384 -4006
rect 4468 -4018 4550 -4006
rect 4966 -4018 5012 -4006
<< via1 >>
rect 2398 610 2468 826
rect 3396 610 3466 826
rect 4392 610 4462 826
rect 988 -4006 1058 -3574
rect 1154 -4008 1224 -3574
rect 1320 -4006 1390 -3572
rect 1486 -4006 1556 -3572
rect 1902 -4006 1972 -3790
rect 2316 -4006 2386 -3572
rect 2482 -4006 2552 -3572
rect 2896 -4006 2966 -3790
rect 3312 -4006 3382 -3572
rect 3478 -4006 3548 -3572
rect 3892 -4006 3962 -3790
rect 4308 -4006 4378 -3572
rect 4474 -4006 4544 -3572
<< metal2 >>
rect 2398 826 2468 836
rect 2398 600 2468 610
rect 3396 826 3466 836
rect 3396 600 3466 610
rect 4392 826 4462 836
rect 4392 600 4462 610
rect 988 -3574 1058 -3564
rect 988 -4016 1058 -4006
rect 1154 -3574 1224 -3564
rect 1154 -4018 1224 -4008
rect 1320 -3572 1390 -3562
rect 1320 -4016 1390 -4006
rect 1486 -3572 1556 -3562
rect 2316 -3572 2386 -3562
rect 1486 -4016 1556 -4006
rect 1902 -3790 1972 -3780
rect 1902 -4016 1972 -4006
rect 2316 -4016 2386 -4006
rect 2482 -3572 2552 -3562
rect 3312 -3572 3382 -3562
rect 2482 -4016 2552 -4006
rect 2896 -3790 2966 -3780
rect 2896 -4016 2966 -4006
rect 3312 -4016 3382 -4006
rect 3478 -3572 3548 -3562
rect 4308 -3572 4378 -3562
rect 3478 -4016 3548 -4006
rect 3892 -3790 3962 -3780
rect 3892 -4016 3962 -4006
rect 4308 -4016 4378 -4006
rect 4474 -3572 4544 -3562
rect 4474 -4016 4544 -4006
<< via2 >>
rect 2398 610 2468 826
rect 3396 610 3466 826
rect 4392 610 4462 826
rect 988 -4006 1058 -3574
rect 1154 -4008 1224 -3574
rect 1320 -4006 1390 -3572
rect 1486 -4006 1556 -3572
rect 1902 -4006 1972 -3790
rect 2316 -4006 2386 -3572
rect 2482 -4006 2552 -3572
rect 2896 -4006 2966 -3790
rect 3312 -4006 3382 -3572
rect 3478 -4006 3548 -3572
rect 3892 -4006 3962 -3790
rect 4308 -4006 4378 -3572
rect 4474 -4006 4544 -3572
<< metal3 >>
rect 2388 826 2478 831
rect 2388 655 2398 826
rect 1892 610 2398 655
rect 2468 655 2478 826
rect 3386 826 3476 831
rect 3386 655 3396 826
rect 2468 610 2479 655
rect 1892 565 2479 610
rect 2886 610 3396 655
rect 3466 655 3476 826
rect 4382 826 4472 832
rect 3466 610 3477 655
rect 4382 654 4392 826
rect 2886 565 3477 610
rect 3883 610 4392 654
rect 4462 610 4472 826
rect 3883 565 4472 610
rect 978 -3574 1068 -3569
rect 978 -4006 988 -3574
rect 1058 -4006 1068 -3574
rect 978 -4011 1068 -4006
rect 1144 -3574 1234 -3569
rect 1144 -4008 1154 -3574
rect 1224 -4008 1234 -3574
rect 1144 -4013 1234 -4008
rect 1310 -3572 1400 -3567
rect 1310 -4006 1320 -3572
rect 1390 -4006 1400 -3572
rect 1310 -4011 1400 -4006
rect 1476 -3572 1566 -3567
rect 1476 -4006 1486 -3572
rect 1556 -4006 1566 -3572
rect 1476 -4011 1566 -4006
rect 1892 -3790 1982 565
rect 1892 -4006 1902 -3790
rect 1972 -4006 1982 -3790
rect 1892 -4011 1982 -4006
rect 2306 -3572 2396 -3567
rect 2306 -4006 2316 -3572
rect 2386 -4006 2396 -3572
rect 2306 -4011 2396 -4006
rect 2472 -3572 2562 -3567
rect 2472 -4006 2482 -3572
rect 2552 -4006 2562 -3572
rect 2472 -4011 2562 -4006
rect 2886 -3790 2976 565
rect 2886 -4006 2896 -3790
rect 2966 -4006 2976 -3790
rect 2886 -4011 2976 -4006
rect 3302 -3572 3392 -3567
rect 3302 -4006 3312 -3572
rect 3382 -4006 3392 -3572
rect 3302 -4011 3392 -4006
rect 3468 -3572 3558 -3567
rect 3468 -4006 3478 -3572
rect 3548 -4006 3558 -3572
rect 3883 -3700 3972 565
rect 3468 -4011 3558 -4006
rect 3882 -3790 3972 -3700
rect 3882 -4006 3892 -3790
rect 3962 -4006 3972 -3790
rect 3882 -4011 3972 -4006
rect 4298 -3572 4388 -3567
rect 4298 -4006 4308 -3572
rect 4378 -4006 4388 -3572
rect 4298 -4011 4388 -4006
rect 4464 -3572 4554 -3567
rect 4464 -4006 4474 -3572
rect 4544 -4006 4554 -3572
rect 4464 -4011 4554 -4006
use sky130_fd_pr__res_high_po_0p35_CN8CXG  sky130_fd_pr__res_high_po_0p35_CN8CXG_0
timestamp 1716574166
transform 1 0 2766 0 1 -1590
box -2276 -2582 2276 2582
<< labels >>
flabel metal3 978 -4010 1068 -3920 0 FreeSans 800 270 0 0 gnd
flabel metal3 1144 -4012 1234 -3922 0 FreeSans 800 270 0 0 vdd
flabel metal3 4382 742 4472 832 0 FreeSans 800 270 0 0 vdac
flabel metal3 1310 -4010 1400 -3920 0 FreeSans 800 90 0 0 i_x8[1]
flabel metal3 1476 -4010 1566 -3920 0 FreeSans 800 90 0 0 i_x8[0]
flabel metal3 2306 -4010 2396 -3920 0 FreeSans 800 90 0 0 i_x4[1]
flabel metal3 2472 -4010 2562 -3920 0 FreeSans 800 90 0 0 i_x4[0]
flabel metal3 3302 -4010 3392 -3920 0 FreeSans 800 90 0 0 i_x2[1]
flabel metal3 3468 -4010 3558 -3920 0 FreeSans 800 90 0 0 i_x2[0]
flabel metal3 4298 -4010 4388 -3920 0 FreeSans 800 90 0 0 i_x1[1]
flabel metal3 4464 -4010 4554 -3920 0 FreeSans 800 90 0 0 i_x1[0]
<< end >>
