magic
tech sky130A
magscale 1 2
timestamp 1716574166
<< pwell >>
rect -2276 -2582 2276 2582
<< psubdiff >>
rect -2240 2512 -2144 2546
rect 2144 2512 2240 2546
rect -2240 2450 -2206 2512
rect 2206 2450 2240 2512
rect -2240 -2512 -2206 -2450
rect 2206 -2512 2240 -2450
rect -2240 -2546 -2144 -2512
rect 2144 -2546 2240 -2512
<< psubdiffcont >>
rect -2144 2512 2144 2546
rect -2240 -2450 -2206 2450
rect 2206 -2450 2240 2450
rect -2144 -2546 2144 -2512
<< xpolycontact >>
rect -2110 1984 -2040 2416
rect -2110 -2416 -2040 -1984
rect -1944 1984 -1874 2416
rect -1944 -2416 -1874 -1984
rect -1778 1984 -1708 2416
rect -1778 -2416 -1708 -1984
rect -1612 1984 -1542 2416
rect -1612 -2416 -1542 -1984
rect -1446 1984 -1376 2416
rect -1446 -2416 -1376 -1984
rect -1280 1984 -1210 2416
rect -1280 -2416 -1210 -1984
rect -1114 1984 -1044 2416
rect -1114 -2416 -1044 -1984
rect -948 1984 -878 2416
rect -948 -2416 -878 -1984
rect -782 1984 -712 2416
rect -782 -2416 -712 -1984
rect -616 1984 -546 2416
rect -616 -2416 -546 -1984
rect -450 1984 -380 2416
rect -450 -2416 -380 -1984
rect -284 1984 -214 2416
rect -284 -2416 -214 -1984
rect -118 1984 -48 2416
rect -118 -2416 -48 -1984
rect 48 1984 118 2416
rect 48 -2416 118 -1984
rect 214 1984 284 2416
rect 214 -2416 284 -1984
rect 380 1984 450 2416
rect 380 -2416 450 -1984
rect 546 1984 616 2416
rect 546 -2416 616 -1984
rect 712 1984 782 2416
rect 712 -2416 782 -1984
rect 878 1984 948 2416
rect 878 -2416 948 -1984
rect 1044 1984 1114 2416
rect 1044 -2416 1114 -1984
rect 1210 1984 1280 2416
rect 1210 -2416 1280 -1984
rect 1376 1984 1446 2416
rect 1376 -2416 1446 -1984
rect 1542 1984 1612 2416
rect 1542 -2416 1612 -1984
rect 1708 1984 1778 2416
rect 1708 -2416 1778 -1984
rect 1874 1984 1944 2416
rect 1874 -2416 1944 -1984
rect 2040 1984 2110 2416
rect 2040 -2416 2110 -1984
<< ppolyres >>
rect -2110 -1984 -2040 1984
rect -1944 -1984 -1874 1984
rect -1778 -1984 -1708 1984
rect -1612 -1984 -1542 1984
rect -1446 -1984 -1376 1984
rect -1280 -1984 -1210 1984
rect -1114 -1984 -1044 1984
rect -948 -1984 -878 1984
rect -782 -1984 -712 1984
rect -616 -1984 -546 1984
rect -450 -1984 -380 1984
rect -284 -1984 -214 1984
rect -118 -1984 -48 1984
rect 48 -1984 118 1984
rect 214 -1984 284 1984
rect 380 -1984 450 1984
rect 546 -1984 616 1984
rect 712 -1984 782 1984
rect 878 -1984 948 1984
rect 1044 -1984 1114 1984
rect 1210 -1984 1280 1984
rect 1376 -1984 1446 1984
rect 1542 -1984 1612 1984
rect 1708 -1984 1778 1984
rect 1874 -1984 1944 1984
rect 2040 -1984 2110 1984
<< locali >>
rect -2240 2512 -2144 2546
rect 2144 2512 2240 2546
rect -2240 2450 -2206 2512
rect 2206 2450 2240 2512
rect -2240 -2512 -2206 -2450
rect 2206 -2512 2240 -2450
rect -2240 -2546 -2144 -2512
rect 2144 -2546 2240 -2512
<< viali >>
rect -2094 2001 -2056 2398
rect -1928 2001 -1890 2398
rect -1762 2001 -1724 2398
rect -1596 2001 -1558 2398
rect -1430 2001 -1392 2398
rect -1264 2001 -1226 2398
rect -1098 2001 -1060 2398
rect -932 2001 -894 2398
rect -766 2001 -728 2398
rect -600 2001 -562 2398
rect -434 2001 -396 2398
rect -268 2001 -230 2398
rect -102 2001 -64 2398
rect 64 2001 102 2398
rect 230 2001 268 2398
rect 396 2001 434 2398
rect 562 2001 600 2398
rect 728 2001 766 2398
rect 894 2001 932 2398
rect 1060 2001 1098 2398
rect 1226 2001 1264 2398
rect 1392 2001 1430 2398
rect 1558 2001 1596 2398
rect 1724 2001 1762 2398
rect 1890 2001 1928 2398
rect 2056 2001 2094 2398
rect -2094 -2398 -2056 -2001
rect -1928 -2398 -1890 -2001
rect -1762 -2398 -1724 -2001
rect -1596 -2398 -1558 -2001
rect -1430 -2398 -1392 -2001
rect -1264 -2398 -1226 -2001
rect -1098 -2398 -1060 -2001
rect -932 -2398 -894 -2001
rect -766 -2398 -728 -2001
rect -600 -2398 -562 -2001
rect -434 -2398 -396 -2001
rect -268 -2398 -230 -2001
rect -102 -2398 -64 -2001
rect 64 -2398 102 -2001
rect 230 -2398 268 -2001
rect 396 -2398 434 -2001
rect 562 -2398 600 -2001
rect 728 -2398 766 -2001
rect 894 -2398 932 -2001
rect 1060 -2398 1098 -2001
rect 1226 -2398 1264 -2001
rect 1392 -2398 1430 -2001
rect 1558 -2398 1596 -2001
rect 1724 -2398 1762 -2001
rect 1890 -2398 1928 -2001
rect 2056 -2398 2094 -2001
<< metal1 >>
rect -2100 2398 -2050 2410
rect -2100 2001 -2094 2398
rect -2056 2001 -2050 2398
rect -2100 1989 -2050 2001
rect -1934 2398 -1884 2410
rect -1934 2001 -1928 2398
rect -1890 2001 -1884 2398
rect -1934 1989 -1884 2001
rect -1768 2398 -1718 2410
rect -1768 2001 -1762 2398
rect -1724 2001 -1718 2398
rect -1768 1989 -1718 2001
rect -1602 2398 -1552 2410
rect -1602 2001 -1596 2398
rect -1558 2001 -1552 2398
rect -1602 1989 -1552 2001
rect -1436 2398 -1386 2410
rect -1436 2001 -1430 2398
rect -1392 2001 -1386 2398
rect -1436 1989 -1386 2001
rect -1270 2398 -1220 2410
rect -1270 2001 -1264 2398
rect -1226 2001 -1220 2398
rect -1270 1989 -1220 2001
rect -1104 2398 -1054 2410
rect -1104 2001 -1098 2398
rect -1060 2001 -1054 2398
rect -1104 1989 -1054 2001
rect -938 2398 -888 2410
rect -938 2001 -932 2398
rect -894 2001 -888 2398
rect -938 1989 -888 2001
rect -772 2398 -722 2410
rect -772 2001 -766 2398
rect -728 2001 -722 2398
rect -772 1989 -722 2001
rect -606 2398 -556 2410
rect -606 2001 -600 2398
rect -562 2001 -556 2398
rect -606 1989 -556 2001
rect -440 2398 -390 2410
rect -440 2001 -434 2398
rect -396 2001 -390 2398
rect -440 1989 -390 2001
rect -274 2398 -224 2410
rect -274 2001 -268 2398
rect -230 2001 -224 2398
rect -274 1989 -224 2001
rect -108 2398 -58 2410
rect -108 2001 -102 2398
rect -64 2001 -58 2398
rect -108 1989 -58 2001
rect 58 2398 108 2410
rect 58 2001 64 2398
rect 102 2001 108 2398
rect 58 1989 108 2001
rect 224 2398 274 2410
rect 224 2001 230 2398
rect 268 2001 274 2398
rect 224 1989 274 2001
rect 390 2398 440 2410
rect 390 2001 396 2398
rect 434 2001 440 2398
rect 390 1989 440 2001
rect 556 2398 606 2410
rect 556 2001 562 2398
rect 600 2001 606 2398
rect 556 1989 606 2001
rect 722 2398 772 2410
rect 722 2001 728 2398
rect 766 2001 772 2398
rect 722 1989 772 2001
rect 888 2398 938 2410
rect 888 2001 894 2398
rect 932 2001 938 2398
rect 888 1989 938 2001
rect 1054 2398 1104 2410
rect 1054 2001 1060 2398
rect 1098 2001 1104 2398
rect 1054 1989 1104 2001
rect 1220 2398 1270 2410
rect 1220 2001 1226 2398
rect 1264 2001 1270 2398
rect 1220 1989 1270 2001
rect 1386 2398 1436 2410
rect 1386 2001 1392 2398
rect 1430 2001 1436 2398
rect 1386 1989 1436 2001
rect 1552 2398 1602 2410
rect 1552 2001 1558 2398
rect 1596 2001 1602 2398
rect 1552 1989 1602 2001
rect 1718 2398 1768 2410
rect 1718 2001 1724 2398
rect 1762 2001 1768 2398
rect 1718 1989 1768 2001
rect 1884 2398 1934 2410
rect 1884 2001 1890 2398
rect 1928 2001 1934 2398
rect 1884 1989 1934 2001
rect 2050 2398 2100 2410
rect 2050 2001 2056 2398
rect 2094 2001 2100 2398
rect 2050 1989 2100 2001
rect -2100 -2001 -2050 -1989
rect -2100 -2398 -2094 -2001
rect -2056 -2398 -2050 -2001
rect -2100 -2410 -2050 -2398
rect -1934 -2001 -1884 -1989
rect -1934 -2398 -1928 -2001
rect -1890 -2398 -1884 -2001
rect -1934 -2410 -1884 -2398
rect -1768 -2001 -1718 -1989
rect -1768 -2398 -1762 -2001
rect -1724 -2398 -1718 -2001
rect -1768 -2410 -1718 -2398
rect -1602 -2001 -1552 -1989
rect -1602 -2398 -1596 -2001
rect -1558 -2398 -1552 -2001
rect -1602 -2410 -1552 -2398
rect -1436 -2001 -1386 -1989
rect -1436 -2398 -1430 -2001
rect -1392 -2398 -1386 -2001
rect -1436 -2410 -1386 -2398
rect -1270 -2001 -1220 -1989
rect -1270 -2398 -1264 -2001
rect -1226 -2398 -1220 -2001
rect -1270 -2410 -1220 -2398
rect -1104 -2001 -1054 -1989
rect -1104 -2398 -1098 -2001
rect -1060 -2398 -1054 -2001
rect -1104 -2410 -1054 -2398
rect -938 -2001 -888 -1989
rect -938 -2398 -932 -2001
rect -894 -2398 -888 -2001
rect -938 -2410 -888 -2398
rect -772 -2001 -722 -1989
rect -772 -2398 -766 -2001
rect -728 -2398 -722 -2001
rect -772 -2410 -722 -2398
rect -606 -2001 -556 -1989
rect -606 -2398 -600 -2001
rect -562 -2398 -556 -2001
rect -606 -2410 -556 -2398
rect -440 -2001 -390 -1989
rect -440 -2398 -434 -2001
rect -396 -2398 -390 -2001
rect -440 -2410 -390 -2398
rect -274 -2001 -224 -1989
rect -274 -2398 -268 -2001
rect -230 -2398 -224 -2001
rect -274 -2410 -224 -2398
rect -108 -2001 -58 -1989
rect -108 -2398 -102 -2001
rect -64 -2398 -58 -2001
rect -108 -2410 -58 -2398
rect 58 -2001 108 -1989
rect 58 -2398 64 -2001
rect 102 -2398 108 -2001
rect 58 -2410 108 -2398
rect 224 -2001 274 -1989
rect 224 -2398 230 -2001
rect 268 -2398 274 -2001
rect 224 -2410 274 -2398
rect 390 -2001 440 -1989
rect 390 -2398 396 -2001
rect 434 -2398 440 -2001
rect 390 -2410 440 -2398
rect 556 -2001 606 -1989
rect 556 -2398 562 -2001
rect 600 -2398 606 -2001
rect 556 -2410 606 -2398
rect 722 -2001 772 -1989
rect 722 -2398 728 -2001
rect 766 -2398 772 -2001
rect 722 -2410 772 -2398
rect 888 -2001 938 -1989
rect 888 -2398 894 -2001
rect 932 -2398 938 -2001
rect 888 -2410 938 -2398
rect 1054 -2001 1104 -1989
rect 1054 -2398 1060 -2001
rect 1098 -2398 1104 -2001
rect 1054 -2410 1104 -2398
rect 1220 -2001 1270 -1989
rect 1220 -2398 1226 -2001
rect 1264 -2398 1270 -2001
rect 1220 -2410 1270 -2398
rect 1386 -2001 1436 -1989
rect 1386 -2398 1392 -2001
rect 1430 -2398 1436 -2001
rect 1386 -2410 1436 -2398
rect 1552 -2001 1602 -1989
rect 1552 -2398 1558 -2001
rect 1596 -2398 1602 -2001
rect 1552 -2410 1602 -2398
rect 1718 -2001 1768 -1989
rect 1718 -2398 1724 -2001
rect 1762 -2398 1768 -2001
rect 1718 -2410 1768 -2398
rect 1884 -2001 1934 -1989
rect 1884 -2398 1890 -2001
rect 1928 -2398 1934 -2001
rect 1884 -2410 1934 -2398
rect 2050 -2001 2100 -1989
rect 2050 -2398 2056 -2001
rect 2094 -2398 2100 -2001
rect 2050 -2410 2100 -2398
<< properties >>
string FIXED_BBOX -2223 -2529 2223 2529
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 20 m 1 nx 26 wmin 0.350 lmin 0.50 rho 319.8 val 19.387k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
